ABS_REG_CFG_MAIN_CLKS, 32'h0012_0023
ABS_REG_DAC_WORK     , 32'd0012_0023
